
module IFlipFlop(iff_in, iff_out);

input iff_in;
output iff_out;

endmodule
